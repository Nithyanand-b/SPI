import uvm_pkg::*;

`include "uvm_macros.svh"
`include "dut/spi_interface.sv"
`include "dut/dut.sv"
`include "dut/spi_config.sv"
`include "testbench/transaction.sv"
`include "testbench/sequences.sv"
`include "testbench/driver.sv"
`include "testbench/monitor.sv"
`include "testbench/scoreboard.sv"
`include "testbench/agent.sv"
`include "testbench/env.sv"
`include "testbench/test.sv"